module capas

fn context_test(){
	mut ctx := 
}