module main

import linklancien.capas

fn main(){}